library ieee;
use ieee.std_logic_1164.all;
entity NOR1BIT is
    Port ( A : in  STD_LOGIC;
 B : in  STD_LOGIC;
 C : out  STD_LOGIC);
end NOR1BIT;
architecture Behavioral of NOR1BIT is
begin
C<= A NOR B;
end�Behavioral;